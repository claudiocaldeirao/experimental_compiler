BEGIN
    x = 5;
    y = x + 2;
    z = y;
    PRINT z;
END
