BEGIN
    x = 5;
    y = x + 2;
    z = y;
END
